

module bypass (
    ports
);
    
endmodule



