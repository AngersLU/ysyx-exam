//write back

//`include "defines.v"

// module wbu (
//     input wire clk,
//     input wire rst,

//     input reg[`RegAddrBus] wb_w_rd_addr,
//     input reg              wb_w_reg_e,
//     input reg[`RegBus]     wb_w_data

// );

//     regfiel regfile0(.clk(clk),
//                      .rst(rst),
//                      .we(wb_w_reg_e),
//                      .waddr(wb_w_rd_addr),
//                      .re1(),
//                      .raddr1(),
//                      .rdata1());

// endmodule
