
// `timescale 1ns/1ns
// module bypass (
//     po
// );
    
// endmodule



