module ysyx_2022040010_add (
    input wire[63:0] add_src1,
    input wire[63:0] add_src2,
    input wire[x:0]  add_op,

    output reg[63:0] add_result
);
    TODO:
endmodule